library IEEE;
use IEEE.std_logic_1164.all;

package alphabet is
    type alphabet is array (0 to 25) of std_logic_vector (7 downto 0); 
end package alphabet;
